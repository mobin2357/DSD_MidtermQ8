library verilog;
use verilog.vl_types.all;
entity Q8TB is
end Q8TB;
